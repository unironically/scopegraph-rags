grammar statix_translate:to_silver;

--------------------------------------------------

aspect production label
top::Label ::= label::String
{}