grammar statix_translate:lang:analysis;

imports statix_translate:lang:abstractsyntax;