grammar regex_noimports:driver;

imports regex_noimports:resolution;

function main
IO<Integer> ::= largs::[String]
{
  return do {
    return 0;
  };
}