grammar statix_translate:translation;

--------------------------------------------------

fun okNameGen String ::= 
  = "ok_" ++ toString(genInt());