grammar statix_translate:to_ocaml;

imports statix_translate:to_ag;
imports statix_translate:lang:abstractsyntax;