grammar lmr1:lmr:nameanalysis1;

imports syntax:lmr1:lmr:abstractsyntax;
imports sg_lib1:src;