grammar lm_semantics_5:nameanalysis;

imports lm_syntax_1:lang:abstractsyntax;
imports sg_lib;