grammar statix_translate:to_ag;

imports statix_translate:lang:abstractsyntax;
imports statix_translate:lang:analysis;