grammar statix_translate:to_silver;

imports statix_translate:to_ag;
imports statix_translate:lang:abstractsyntax;