grammar statix_translate:translation;

nonterminal Equation;