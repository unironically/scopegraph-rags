grammar lm_semantics_1:nameanalysis;

imports lm_syntax_1:lang:abstractsyntax;