grammar statix_translate:to_silver;

imports statix_translate:lang:abstractsyntax;
imports statix_translate:lang:analysis;