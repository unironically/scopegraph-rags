grammar lmr0:lmr:nameanalysis;

imports syntax:lmr0:lmr:abstractsyntax;
imports sg_lib:src;