grammar lmr0:lmr:nameanalysis1;

imports syntax:lmr0:lmr:abstractsyntax;
imports sg_lib:src;