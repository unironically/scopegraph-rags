grammar statix_translate:translation_two;

imports statix_translate:lang:abstractsyntax;