grammar statix_translate:to_ag;

--------------------------------------------------

aspect production label
top::Label ::= label::String
{}