grammar statix_translate:translation;

imports statix_translate:lang:abstractsyntax;