grammar statix_translate:to_ocaml;

imports statix_translate:to_ag;