imports statix_translate:lang:abstractsyntax;