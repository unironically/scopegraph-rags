grammar lm_semantics_4:nameanalysis;

imports lm_syntax_2:lang:abstractsyntax;
imports sg_lib;