grammar regex_noimports:driver;
imports lmr:lang;

function main
IO<Integer> ::= largs::[String]
{
  return do {
    return 0;
  };
}