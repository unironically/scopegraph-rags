grammar LM;


{-
 - DFA for VarRefs.
 -}
global dfaVarRef::DFA = 
  let sink::State = sinkState() in
  let final::State = state(sink, sink, sink, sink, true) in
  let impState::State = state(final, sink, sink, sink, false) in
  let start::State = state(final, sink, impState, start, false) in
    dfa (start)
  end end end end;

{-
 - DFA for qualified VarRefs.
 -}
global dfaVar::DFA = 
  let final::State = state(sink, sink, sink, sink, true) in
  let start::State = state(final, sink, sink, sink, false) in
    dfa (start)
  end end;

{-
 - DFA for ModRefs.
 -}
global dfaModRef::DFA = 
  let sink::State = sinkState() in
  let final::State = state(sink, sink, sink, sink, true) in
  let impState::State = state(sink, final, sink, sink, false) in
  let start::State = state(sink, final, impState, start, false) in
    dfa (start)
  end end end end;

{-
 - DFA for qualified ModRefs.
 -}
global dfaMod::DFA = 
  let final::State = state(sink, sink, sink, sink, true) in
  let start::State = state(sink, final, sink, sink, false) in
    dfa (start)
  end end;


synthesized attribute findReachable::([Res] ::= String Either<ModRef, VarRef> [Label] Scope);


nonterminal DFA with findReachable;

{-
 - DFA.
 - We only need to hold the start state, as each state knows whether it is final, and there should
 - be a path from the start state to any other state in the DFA.
 -}
abstract production dfa
top::DFA ::=
  start::State
{
  top.findReachable = start.findReachable;
}


nonterminal State with findReachable;

{-
 - Regular (non-sink) state in a DFA.
 - We continue traversal, and also take into account the current scope as a possible resolution
 - if the state is final.
 -}
abstract production state
top::State ::=
  var::State
  mod::State
  imp::State
  lex::State
  isFinal::Boolean
{
  top.findReachable = 
    \lookup::String
     ref::Either<ModRef, VarRef>
     currentPath::[Label]
     currentScope::Scope ->
    
      let varRes::[Res] = if ref.isLeft then [] 
                          else concat(map((var.findReachable(lookup, ref, labelVar()::currentPath, resolvingImp, _)), currentScope.vars)) in
      
      let modRes::[Res] = if ref.isRight then [] 
                          else concat(map((mods.findReachable(lookup, ref, labelMod()::currentPath, resolvingImp, _)), currentScope.mods)) in


      {- `valid` is all of the known reachable import resolutions whose origin is NOT
         equal to the ModRef which we are currently looking up. Then using `valid` in
         the assignment to `imps` below means that the resolution of an import can NOT
         use the IMP edge introduced by itself on a previous iteration of the circ attr. -}
      let valid::[Res] = filter ((\r::Res -> ref.isLeft && r != ref.fromLeft.fromRef),
                                 currentScope.impsReachable) in
      let imps::[Scope] = if ref.isRight then map((.resolvedScope), valid)
                          else scope.imps in
      let impRes::[Res] = concat(map((imps.findReachable(lookup, ref, labelImp()::currentPath, resolvingImp, _)), imps)) in


      let lexRes::[Res] = concat(map((lexs.findReachable(lookup, ref, labelLex()::currentPath, resolvingImp, _)), currentScope.lexs)) in

      let contRes::[Res] = varRef ++ modRes ++ impRes ++ lexRes in

        case currentScope of
        | scopeDatum(d) -> if !isFinal || d.id != lookup then contRes 
                           else if ref.isLeft then impRes(left(ref), currentScope, currentPath) :: contRes
                           else varRes(right(ref), currentScope, currentPath) :: contRes 
        | _ -> contRes -- ignore scopes that do not have data
        end

      end end end end end end end;
}

{-
 - Sink state in a DFA. 
 - Cannot use the current scope in a resolution, and cannot transition.
 -}
abstract production sinkState
top::State ::=
{
  top.findReachable = 
    \lookup::String 
     ref::Either<ModRef, VarRef> 
     currentPath::[Label] 
     currentScope::Scope -> 
      [];
}
