grammar src_old;