grammar lm_semantics_2:nameanalysis;

imports lm_syntax_2:lang:abstractsyntax;