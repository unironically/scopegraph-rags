grammar lmr1:lmr:nameanalysis5;

imports syntax:lmr1:lmr:abstractsyntax;

import silver:langutil; -- for location.unparse

--------------------------------------------------

monoid attribute ok::Boolean with true, &&;

inherited attribute scope::Decorated Scope;

synthesized attribute VAR_s::[Decorated Scope];
synthesized attribute LEX_s::[Decorated Scope];
synthesized attribute MOD_s::[Decorated Scope];
synthesized attribute IMP_s::[Decorated Scope];

synthesized attribute type::Type;

synthesized attribute module::Maybe<Decorated Scope>;

--------------------------------------------------

attribute ok occurs on Main;

propagate ok on Main;

aspect production program
top::Main ::= ds::Decls
{
  production attribute globScope::Scope = scopeNoData();
  globScope.lex = [];
  globScope.var = [];
  globScope.mod = [];
  globScope.imp = [];

  ds.scope = globScope;
}

--------------------------------------------------

attribute ok, scope, VAR_s, MOD_s occurs on Decls;

propagate ok on Decls;

aspect production declsCons
top::Decls ::= d::Decl ds::Decls
{
  production attribute seqScope::Scope = scopeNoData();
  seqScope.lex = [top.scope];
  seqScope.var = d.VAR_s;
  seqScope.mod = d.MOD_s;
  seqScope.imp = d.IMP_s;

  d.scope = top.scope;
  ds.scope = seqScope;

  top.VAR_s = d.VAR_s ++ ds.VAR_s;
  top.MOD_s = d.MOD_s ++ ds.MOD_s;
}

aspect production declsNil
top::Decls ::=
{
  top.VAR_s = [];
  top.MOD_s = [];
}

--------------------------------------------------

attribute scope occurs on Decl;

attribute VAR_s occurs on Decl;
attribute MOD_s occurs on Decl;
attribute IMP_s occurs on Decl;

attribute ok occurs on Decl;
propagate ok on Decl;

aspect production declModule
top::Decl ::= id::String ds::Decls
{
  production attribute modScope::Scope = scopeMod(id);
  modScope.lex = [top.scope];
  modScope.var = ds.VAR_s;
  modScope.mod = ds.MOD_s;
  modScope.imp = [];

  top.VAR_s = [];
  top.MOD_s = [modScope];
  top.IMP_s = [];

  -- lmr1: variable references should not be able to resolve using the decl
  -- nodes that are defined by ds.VAR_s or ds.MOD_s, breaks forward referencing.
  -- so introduce a different scope to pass down to ds that does not have these

  production attribute lookupScope::Scope = scopeNoData();
  lookupScope.lex = [top.scope];
  lookupScope.var = [];
  lookupScope.mod = [];
  lookupScope.imp = [];

  ds.scope = lookupScope;
}

aspect production declImport
top::Decl ::= r::ModRef
{
  r.scope = top.scope;

  top.VAR_s = [];
  top.MOD_s = [];
  top.IMP_s = case r.module of
              | just(s) -> [s]
              | _ -> []
              end;
}

aspect production declDef
top::Decl ::= b::ParBind
{
  b.scope = top.scope;

  top.VAR_s = b.VAR_s;
  top.MOD_s = [];
  top.IMP_s = [];
}

--------------------------------------------------

attribute scope occurs on Expr;

attribute type occurs on Expr;

attribute ok occurs on Expr;
propagate ok on Expr;

aspect production exprInt
top::Expr ::= i::Integer
{
  top.type = tInt();
}

aspect production exprTrue
top::Expr ::=
{
  top.type= tBool();
}

aspect production exprFalse
top::Expr ::=
{
  top.type= tBool();
}

aspect production exprVar
top::Expr ::= r::VarRef
{
  propagate scope;

  top.type = r.type;
}

aspect production exprAdd
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tInt(), tInt() -> (true, tInt())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprSub
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tInt(), tInt() -> (true, tInt())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprMul
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tInt(), tInt() -> (true, tInt())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprDiv
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tInt(), tInt() -> (true, tInt())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprAnd
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tBool(), tBool() -> (true, tBool())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprOr
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tBool(), tBool() -> (true, tBool())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprEq
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | t1, t2 when t1 == t2 -> (true, tBool())
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprApp
top::Expr ::= e1::Expr e2::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type of
                                   | tFun(t1, t2), t3 when ^t1 == t3 -> (true, ^t2)
                                   | _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprIf
top::Expr ::= e1::Expr e2::Expr e3::Expr
{
  propagate scope;

  local okAndTy::(Boolean, Type) = case e1.type, e2.type, e3.type of
                                   | tBool(), t2, t3 when t2 == t3 -> (true, t2)
                                   | _, _, _ -> (false, tErr())
                                   end;

  top.ok <- okAndTy.1;
  top.type = okAndTy.2;
}

aspect production exprFun
top::Expr ::= d::ArgDecl e::Expr
{
  production attribute bodyScope::Scope = scopeNoData();
  bodyScope.lex = [top.scope];
  bodyScope.var = d.VAR_s;
  bodyScope.mod = [];
  bodyScope.imp = [];

  d.scope = top.scope;
  e.scope = bodyScope;

  top.type = tFun(d.type, e.type);
}

aspect production exprLet
top::Expr ::= bs::SeqBinds e::Expr
{
  production attribute letScope::Decorated Scope = bs.lastScope;

  bs.scope = top.scope;
  e.scope = letScope;

  top.type = e.type;
}

aspect production exprLetRec
top::Expr ::= bs::ParBinds e::Expr
{
  production attribute letScope::Scope = scopeNoData();
  letScope.lex = [top.scope];
  letScope.var = bs.VAR_s;
  letScope.mod = [];
  letScope.imp = [];


  bs.scope = letScope;
  e.scope = letScope;

  top.type = e.type;
}

aspect production exprLetPar
top::Expr ::= bs::ParBinds e::Expr
{
  production attribute letScope::Scope = scopeNoData();
  letScope.lex = [top.scope];
  letScope.var = bs.VAR_s;
  letScope.mod = [];
  letScope.imp = [];

  bs.scope = top.scope;
  e.scope = letScope;

  top.type = e.type;
}

--------------------------------------------------

attribute ok, scope, lastScope occurs on SeqBinds;

propagate ok on SeqBinds;

synthesized attribute lastScope::Decorated Scope;

aspect production seqBindsNil
top::SeqBinds ::=
{
  top.lastScope = top.scope;
}

aspect production seqBindsOne
top::SeqBinds ::= s::SeqBind
{
  production attribute sbScope::Scope = scopeNoData();
  sbScope.lex = [top.scope];
  sbScope.var = s.VAR_s;
  sbScope.mod = [];
  sbScope.imp = [];

  s.scope = top.scope;

  top.lastScope = sbScope;
}

aspect production seqBindsCons
top::SeqBinds ::= s::SeqBind ss::SeqBinds
{
  production attribute sbScope::Scope = scopeNoData();
  sbScope.lex = [top.scope];
  sbScope.var = s.VAR_s;
  sbScope.mod = [];
  sbScope.imp = [];

  s.scope = top.scope;
  ss.scope = sbScope;

  top.lastScope = ss.lastScope;
}

--------------------------------------------------

attribute ok, scope, VAR_s occurs on SeqBind;

propagate ok on SeqBind;

aspect production seqBindUntyped
top::SeqBind ::= id::String e::Expr
{
  production attribute varScope::Scope = scopeVar(id, e.type);
  varScope.lex = [];
  varScope.var = [];
  varScope.mod = [];
  varScope.imp = [];

  e.scope = top.scope;

  top.VAR_s = [varScope];
}

aspect production seqBindTyped
top::SeqBind ::= ty::Type id::String e::Expr
{
  production attribute varScope::Scope = scopeVar(id, ^ty);
  varScope.lex = [];
  varScope.var = [];
  varScope.mod = [];
  varScope.imp = [];

  e.scope = top.scope;

  top.ok <- e.type == ^ty;
  top.VAR_s = [varScope];
}

--------------------------------------------------

attribute ok, scope, VAR_s occurs on ParBinds;

propagate ok, scope on ParBinds;

aspect production parBindsNil
top::ParBinds ::=
{
  top.VAR_s = [];
}

aspect production parBindsCons
top::ParBinds ::= s::ParBind ss::ParBinds
{
  top.VAR_s = s.VAR_s ++ ss.VAR_s;
}

--------------------------------------------------

attribute ok, scope, VAR_s occurs on ParBind;

propagate ok on ParBind;

aspect production parBindUntyped
top::ParBind ::= id::String e::Expr
{
  production attribute varScope::Scope = scopeVar(id, e.type);
  varScope.lex = [];
  varScope.var = [];
  varScope.mod = [];
  varScope.imp = [];

  e.scope = top.scope;

  top.VAR_s = [varScope];
}

aspect production parBindTyped
top::ParBind ::= ty::Type id::String e::Expr
{
  production attribute varScope::Scope = scopeVar(id, ^ty);
  varScope.lex = [];
  varScope.var = [];
  varScope.mod = [];
  varScope.imp = [];

  e.scope = top.scope;

  top.ok <- e.type == ^ty;
  top.VAR_s = [varScope];
}

--------------------------------------------------

attribute ok, scope, type, VAR_s occurs on ArgDecl;

propagate ok on ArgDecl;

aspect production argDecl
top::ArgDecl ::= id::String tyann::Type
{
  production attribute varScope::Scope = scopeVar(id, ^tyann);
  varScope.lex = [];
  varScope.var = [];
  varScope.mod = [];
  varScope.imp = [];

  top.type = ^tyann;
  top.VAR_s = [varScope];
}

--------------------------------------------------

aspect production tFun
top::Type ::= tyann1::Type tyann2::Type
{}

aspect production tInt
top::Type ::=
{}

aspect production tBool
top::Type ::=
{}

aspect production tErr
top::Type ::=
{}

--------------------------------------------------

attribute ok, scope, type occurs on VarRef;

aspect production varRef
top::VarRef ::= x::String
{
  local xvars_::[Decorated Scope] =
    top.scope.resolve(isName(x), varRx(), labelOrd);

  local okAndRes::(Boolean, Type) = 
    if length(xvars_) < 1
    then unsafeTracePrint((false, tErr()), "[✗] " ++ top.location.unparse ++ 
                          ": error: unresolvable variable reference '" ++ x ++ "'\n")
    else if length(xvars_) > 1
    then unsafeTracePrint((false, tErr()), "[✗] " ++ top.location.unparse ++ 
                          ": error: ambiguous variable reference '" ++ x ++ "'\n")
    else case head(xvars_).datum of
         | datumVar(_, ty) -> (true, ^ty)
         | _ -> (false, tErr())
         end;

  top.ok := okAndRes.1;
  top.type = okAndRes.2;
}

--------------------------------------------------

attribute scope, ok, module occurs on ModRef;

aspect production modRef
top::ModRef ::= x::String
{
  local xmods_::[Decorated Scope] =
    top.scope.resolve(isName(x), modRx(), labelOrd);

  local okAndRes::(Boolean, Maybe<Decorated Scope>) = 
    if length(xmods_) < 1
    then unsafeTracePrint((false, nothing()), "[✗] " ++ top.location.unparse ++ 
                          ": error: unresolvable module reference '" ++ x ++ "'\n")
    else if length(xmods_) > 1
    then unsafeTracePrint((false, nothing()), "[✗] " ++ top.location.unparse ++ 
                          ": error: ambiguous module reference '" ++ x ++ "'\n")
    else case head(xmods_).datum of
         | datumMod(_) -> (true, just(head(xmods_)))
         | _ -> (false, nothing())
         end;

  top.ok := okAndRes.1;
  top.module = okAndRes.2;
}