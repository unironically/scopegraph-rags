grammar LM;

collection attribute binds::[(String, String)] with ++, [] root Program;

