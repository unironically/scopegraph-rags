grammar lm_semantics_3:nameanalysis;

imports lm_syntax_2:lang:abstractsyntax;