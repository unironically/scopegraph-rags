grammar LM;

--EVW: this is also declared in LM_Scoping.sv
collection attribute binds::[(String, String)] with ++, [] root Program;

