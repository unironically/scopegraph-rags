../../../statix_translate/silver_ag.sv