grammar lm_semantics_0:nameanalysis;

imports lm_syntax_0:lang:abstractsyntax;
imports sg_lib;