grammar statix_translate:translation;

--------------------------------------------------

synthesized attribute refNamesList::[String] occurs on RefNameList;

aspect production refNameListCons
top::RefNameList ::= name::String names::RefNameList
{
  top.refNamesList = name :: names.refNamesList;
}

aspect production refNameListOne
top::RefNameList ::= name::String
{
  top.refNamesList = [name];
}

--------------------------------------------------

synthesized attribute nameListDefs::[(String, TypeAnn)] occurs on NameList;

aspect production nameListCons
top::NameList ::= name::Name names::NameList
{
  top.nameListDefs = name.nameDef :: names.nameListDefs;
}

aspect production nameListOne
top::NameList ::= name::Name
{
  top.nameListDefs = [name.nameDef];
}


synthesized attribute nameDef::(String, TypeAnn) occurs on Name;

aspect production nameSyn
top::Name ::= name::String ty::TypeAnn
{
  top.nameDef = (name, ^ty);
}

aspect production nameInh
top::Name ::= name::String ty::TypeAnn
{
  top.nameDef = (name, ^ty);
}

aspect production nameRet
top::Name ::= name::String ty::TypeAnn
{
  top.nameDef = (name, ^ty);
}

aspect production nameUntagged
top::Name ::= name::String ty::TypeAnn
{
  top.nameDef = (name, ^ty);
}